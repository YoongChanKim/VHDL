LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY TB_BINARYCOMPARATOR IS
END TB_BINARYCOMPARATOR;
ARCHITECTURE HB OF TB_BINARYCOMPARATOR IS
COMPONENT BINARYCOMPARATOR
PORT (
	A,B : IN BIT;
	G1,G2,G3 : OUT BIT
	);
END COMPONENT;
SIGNAL A : BIT := '0';
SIGNAL B : BIT := '0';

SIGNAL G1 : BIT := '0';
SIGNAL G2 : BIT := '0';
SIGNAL G3 : BIT := '0';

BEGIN 
A <='0', '0' AFTER 100NS, '0' AFTER 200NS, '1' AFTER 300NS, '1' AFTER 400NS;
B <='0', '0' AFTER 100NS, '1' AFTER 200NS, '0' AFTER 300NS, '1' AFTER 400NS;

U_BINARYCOMPARATOR : BINARYCOMPARATOR
PORT MAP (
	A => A,
	B => B,
	
	G1 => G1,
	G2 => G2,
	G3 => G3
);
END HB;
