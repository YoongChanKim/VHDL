--TB_HB_FA.VHD 
LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_HB_EXAMPLE IS
END TB_HB_EXAMPLE;

ARCHITECTURE HB OF TB_HB_EXAMPLE IS
	COMPONENT HB_HA IS
	PORT(
			A,B:IN BIT; 
			Y : OUT BIT
	);
	END COMPONENT;
	
	SIGNAL A,B :BIT:='0';
	SIGNAL Y :BIT:='0';
	
	BEGIN
	A <= '0','0' AFTER 100NS,'0' AFTER 200NS,'1' AFTER 300NS, '1' AFTER 400NS,
	B <= '0','0' AFTER 100NS,'1' AFTER 200NS,'0' AFTER 300NS, '1' AFTER 400NS,
	
	U_HB_EXAMPLE : HB_EXAMPLE 
	PORT MAP(
		A=>A,
		B=>B,
		Y=>Y
	);
	END HB;
	