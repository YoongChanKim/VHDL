ENTITY HB_AND2 IS
PORT(
	A,B : IN BIT;
	X : OUT BIT;
	y : OUT BIT
);

END HB_AND2;

ARCHITECTURE HB OF HB_AND2 IS
BEGIN
	X <= A AND B;
	Y <= A OR B;
	
END HB;