ENTITY BINARYCOMPARATOR IS
PORT(
	A,B : IN BIT;
	G1,G2,G3 : OUT BIT
	);
	END BINARYCOMPARATOR;
	
	ARCHITECTURE HB OF BINARYCOMPARATOR IS
	BEGIN 
	
	G1 <= A AND (NOT B);
	G2 <= A XNOR B;
	G3 <= B AND (NOT A);
	
	END HB;
	
	