LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY TB_HB_SEG_DECODER IS
END TB_HB_SEG_DECODER; 
ARCHITECTURE HB OF TB_HB_SEG_DECODER IS 
COMPONENT HB_SEG_DECODER
 PORT ( 
	BCD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 a, b, c, d, e, f, g : OUT STD_LOGIC 
); 
END COMPONENT; 
SIGNAL 
	BCD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000"; 
	SIGNAL A, B, C, D : STD_LOGIC; 
	SIGNAL E, F, G : STD_LOGIC; 
BEGIN
 BCD <= "0000", "0001" AFTER 100NS, "0010" AFTER 200NS, "0011" AFTER 300NS, "0100" AFTER 
               400NS, "0101" AFTER 500NS, "0110" AFTER 600NS, "0111" AFTER 700NS, "1000" AFTER 
               800NS, "1001" AFTER 900NS; 
U_HB_SEG_DECODER : HB_SEG_DECODER 
PORT MAP ( 
           BCD => BCD, A => A, B => B, C => C, D => D, E => E, F => F, G => G 
);
 END HB; 	
