
ENTITY HB_EXAMPLE IS
PORT(
	A,B : IN BIT;
	Y : OUT BIT 
);
END EXAMPLE;

ARCHITECTURE HB OF HB_EXAMPLE IS
	COMPONENT HB_HA IS
	PORT(
			A,B:IN BIT; 
			Y : OUT BIT
	);
	END COMPONENT;
	SIGNAL X1,X2,X3:BIT;
	
	BEGIN
	PORT MAP(
		X1 <= A NAND B;
		X2 <= A NAND X1;
		X3 <= B NAND X2;
		Y  <= X2 NAND X3
		);
		END HB;
		
		